module decoder_2x4_sheffer (input [1:0] a, output [3:0] b);
wire [3:0] nb;

 assign nb[3] = ~(~(a[1] & a[0]) & ~(a[1] & a[0])),
        nb[2] = ~(~(a[1] & ~(a[0] & a[0])) & 
                  ~(a[1] & ~(a[0] & a[0]))),  
        nb[1] = ~(~(~(a[1] & a[1]) & a[0]) & 
                  ~(~(a[1] & a[1]) & a[0])),
        nb[0] = ~(~(~(a[1] & a[1]) & ~(a[0] &
                a[0])) & ~(~(a[1] & a[1]) & ~(a[0] & a[0]))),
         b[3] = ~(nb[3] & nb[3]), 
         b[2] = ~(nb[2] & nb[2]), 
         b[1] = ~(nb[1] & nb[1]), 
         b[0] = ~(nb[0] & nb[0]); 

endmodule